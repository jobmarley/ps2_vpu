
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity vpu_test_simul is
--  Port ( );
end vpu_test_simul;

architecture vpu_test_simul_behavioral of vpu_test_simul is
 component design_4 is
  end component design_4;
begin
design_4_i: component design_4
 ;

end vpu_test_simul_behavioral;
